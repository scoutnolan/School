entity CONVERTER is
  port (B:in bit_vector (3 downto 0);
        E: out bit_vector (3 downto 0));
end CONVERTER;
