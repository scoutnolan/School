configuration STRUCTURAL of TEST_BENCH is
  for CONVERTER_TEST
    for L1 : CONVERTERC 
      use entity CONVERTER(STRUCTURAL);
    end for;
  end for;
end STRUCTURAL;
